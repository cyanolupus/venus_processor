module exec_ldst ();
    
endmodule